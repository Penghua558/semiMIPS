/*
* File Name: idexreg_tb.v
* Function: this is a testbench file for module ID/EX pipeline register.
*/

module idexreg_tb ();
endmodule
